// responsible for returning the 32 bit instruction assosciated with the PC
// will read from a plaintext file that contains the instructions. those instructions will be stored in a related
module programmemory

endmodule